package tp is
--constant numBit : integer := 11;
constant N : integer  := 8;
constant NB : integer := 11;
constant SHAMT : integer := 12;

end tp ;